# ====================================================================
#
#      99685.cdl
#
#      Compact flash interface camera
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2004 Winbond.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      clyu
# Contributors:   clyu
# Date:           2004-8-23
#
#####DESCRIPTIONEND####

cdl_package CYGPKG_DEVS_MEDIA_VIDEO_W99685 {
    display       "w99685 device driver"
    description   "w99685 camera driver for CFI interface"

    requires      CYGPKG_IO
    requires      CYGPKG_IO_W99685
    requires      CYGPKG_ISOINFRA
    requires      CYGINT_ISO_C_TIME_TYPES
    requires      CYGINT_ISO_STRERROR
    requires      CYGINT_ISO_ERRNO
    requires      CYGINT_ISO_ERRNO_CODES
    requires      CYGINT_ISO_MALLOC
    requires      CYGPKG_LINUX_COMPAT
    requires	  CYGPKG_IO_FILEIO

    include_dir   video

	implements    CYGHWR_IO_SDRAM_DEVICE
	compile      -library=libextras.a w99685.c
	
	cdl_option CYGPKG_MEDIA_VIDEO_W99685_FUNCTIONS {
		display "w99685 functions support"
        default_value 1
        	
		compile		w99685CFI.c
    	description "
            w99685 functions support."
    }
    cdl_option CYGDAT_MEDIA_VIDEO_VIDEO0_NAME {
    	display "w99685 device name"
        flavor        data
	    default_value {"\"/dev/video0\""}
        	
    	description "
            This option specifies the name of the w99685 device for the 
            ARM W90N740."
    }
    
	cdl_component CYGPKG_MEDIA_VIDEO_W99685_SENSOR {
        display "sensor"
        default_value 1

        description "
            support which sensor."
		
		
        cdl_option CYGPKG_MEDIA_VIDEO_W99685_SS {
	        display "SumSung sensor support"
        	default_value 1

    	    description "
            SumSung sensor support."
    	}
    	cdl_option CYGPKG_MEDIA_VIDEO_W99685_OV {
	        display "OV sensor support"
        	default_value 0

    	    description "
            OV sensor support."
    	}
    	cdl_option CYGPKG_MEDIA_VIDEO_W99685_HYNIX {
	        display "HYNIX sensor support"
        	default_value 0

    	    description "
            HYNIX sensor support."
    	}
    	cdl_option CYGPKG_MEDIA_VIDEO_W99685_TS {
	        display "ToShiBa sensor support"
        	default_value 0

    	    description "
            ToShiBa sensor support."
    	}
    }
    
	cdl_component CYGPKG_DEVS_MEDIA_VIDEO_W99685_OPTIONS {
        display "W99685 support build options"
        flavor  none
        no_define

        cdl_option CYGPKG_DEVS_MEDIA_VIDEO_W99685_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the networking package.
                These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_MEDIA_VIDEO_W99685_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the networking package. These flags are removed from
                the set of global flags if present."
        }
    }
}

