# ====================================================================
#
#      ser_arm_integrator.cdl
#
#      eCos serial ARM/INTEGRATOR configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      David A Rusling
# Original data:  David A Rusling
# Contributors:	  Philippe Robin
# Date:           November 7, 2000
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_ARM_INTEGRATOR {
    display       "ARM INTEGRATOR serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_ARM_INTEGRATOR

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    description   "
           This option enables the serial device drivers for the
           ARM INTEGRATOR."

    compile       -library=libextras.a   integrator_serial_with_ints.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_arm_integrator.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_INTEGRATOR_SERIAL0 {
	display       "ARM INTEGRATOR serial port 0 driver"
	flavor        bool
	default_value 1
	description   "
        This option includes the serial device driver for the ARM INTEGRATOR 
        port 0."

	cdl_option CYGDAT_IO_SERIAL_ARM_INTEGRATOR_SERIAL0_NAME {
	    display       "Device name for ARM INTEGRATOR serial port 0 driver"
	    flavor        data
	    default_value {"\"/dev/ser0\""}
	    description   "
            This option specifies the name of the serial device for the 
            ARM INTEGRATOR port 0."
	}

	cdl_option CYGNUM_IO_SERIAL_ARM_INTEGRATOR_SERIAL0_BAUD {
	    display       "Baud rate for the ARM INTEGRATOR serial port 0 driver"
	    flavor        data
	    legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
	    		    4800 7200 9600 14400 19200 38400 57600 115200 234000
			   }
	    default_value 38400
	    description   "
            This option specifies the default baud rate (speed) for the 
            ARM INTEGRATOR port 0."
	}

	cdl_option CYGNUM_IO_SERIAL_ARM_INTEGRATOR_SERIAL0_BUFSIZE {
	    display       "Buffer size for the ARM INTEGRATOR serial port 0 driver"
	    flavor        data
	    legal_values  0 to 8192
	    default_value 128
	    description   "
            This option specifies the size of the internal buffers used 
            for the ARM INTEGRATOR port 0."
	}
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_INTEGRATOR_SERIAL1 {
	display       "ARM INTEGRATOR serial port 1 driver"
	flavor        bool
	default_value 1
	description   "
        This option includes the serial device driver for the ARM INTEGRATOR 
        port 1."

	cdl_option CYGDAT_IO_SERIAL_ARM_INTEGRATOR_SERIAL1_NAME {
	    display       "Device name for ARM INTEGRATOR serial port 1 driver"
	    flavor        data
	    default_value {"\"/dev/ser1\""}
	    description   "
            This option specifies the name of the serial device for the 
            ARM INTEGRATOR port 1."
	}

	cdl_option CYGNUM_IO_SERIAL_ARM_INTEGRATOR_SERIAL1_BAUD {
	    display       "Baud rate for the ARM INTEGRATOR serial port 1 driver"
	    flavor        data
	    legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 234000
            }
	    default_value 38400
	    description   "
            This option specifies the default baud rate (speed) for the
            ARM INTEGRATOR port 1."
	}
    }

    cdl_option CYGNUM_IO_SERIAL_ARM_INTEGRATOR_SERIAL1_BUFSIZE {
        display       "Buffer size for the ARM INTEGRATOR serial port 1 driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the ARM INTEGRATOR port 1."
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_INTEGRATOR_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_ARM_INTEGRATOR_SERIAL0

	# The combination of non-FIFO UARTs and no cache means that some 
	# Integrator based systems are too slow to handle the higher baud rates.
        implements CYGINT_IO_SERIAL_TEST_SKIP_57600
	implements CYGINT_IO_SERIAL_TEST_SKIP_115200
	
        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_ARM_INTEGRATOR_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"arminteg\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF ser_arm_integrator.cdl
