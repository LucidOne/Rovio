# ====================================================================
#
#      profile_gprof.cdl
#
#      cpu load measurements
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2002 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Gary Thomas
# Original data:  Gary Thomas
# Contributors:
# Date:           2002-11-14
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_PROFILE_GPROF {
    display       "Gather runtime profile statistics"
    requires      CYGPKG_NET
    requires      CYGPKG_NET_TFTP
    requires      CYGPKG_MEMALLOC   
    requires      { CYGINT_PROFILE_HAL_TIMER != 0 }
    doc           ref/services-profile-gprof.html

    include_dir   cyg/profile
    
    compile profile.c

    description "
        This package enables runtime profiling of an application.
    The actual profile collection must be turned on by the application,
    once it has been initialized.  The data collected is exported via
    a TFTP connection to the target."

    cdl_interface     CYGINT_PROFILE_HAL_TIMER {
        display   "High resolution timer, implemented by platform"
        description "
	  Profiling requires access to a high resolution timer which
          is platform dependent."
    }

    cdl_option CYGNUM_PROFILE_TFTP_PORT {
        display       "Port used by TFTP server for profile data"
        flavor        data
        default_value 0
        description   "
            This option sets the port number to use for the TFTP server
            which exports the profiling data.  A value of 0 will set
            the port to be the IETF standard port of 69/udp."
    }

    cdl_option CYGPKG_PROFILE_TESTS {
        display "Profiling tests"
        flavor  data   
        no_define      
        calculated { "tests/profile.c" }
    }
}

