# ====================================================================
#
#      io.cdl
#
#      eCos IO configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Original data:  gthomas
# Contributors:
# Date:           1999-07-07
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO {
    display       "I/O sub-system"
    doc           ref/io.html
    include_dir   cyg/io
    requires      CYGPKG_ERROR
    description   "
        The eCos system is supplied with a number of different
        device drivers.  This option enables the basic I/O system
        support which is the basis for all drivers."

    compile       -library=libextras.a ioinit.cxx
    compile       iosys.c

 
    cdl_option CYGDBG_IO_INIT {
        display       "Debug I/O sub-system"
        default_value 0
        description   "
            This option enables verbose messages to be displayed on the
            system 'diag' device during I/O system initialization."
   }

   cdl_component CYGPKG_IO_FILE_SUPPORT {
       display    "Basic support for file based I/O"
       active_if  !CYGPKG_IO_FILEIO
       default_value 1       
       description "
           This option control support for simple file I/O primitives. It is only
           present if the FILEIO package is not included."

       compile       io_file.c

       cdl_option CYGPKG_IO_NFILE {
	   display "Number of open files"
	   flavor  data
	   default_value 16
	   description   "
	       This option controls the number of open files."
       }
    }
}
