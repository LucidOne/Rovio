# ====================================================================
#
#      fat.cdl
#
#      FAT Filesystem configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      clyu
# Date:           2003-12-16
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_FS_FAT {
    display        "FAT filesystem"
    doc            ref/fileio.html
    include_dir    ""

    requires       CYGPKG_IO_FILEIO
    requires       CYGPKG_COMPRESS_ZLIB
    requires       CYGINT_ISO_MALLOC

    requires       CYGPKG_ISOINFRA
    requires       CYGPKG_ERROR
    requires       CYGINT_ISO_ERRNO
    requires       CYGINT_ISO_ERRNO_CODES
    requires       CYGPKG_IO_FILEIO_INODE
    requires       CYGPKG_LINUX_COMPAT
    requires       CYGPKG_CRC

    implements     CYGINT_IO_FILEIO_FS      

    compile        blockio.c  drives.c fat16.c readdir.c \
				   creat.c fat32.c lfn.c readwrit.c \
				   attrib.c  mount.c request.c \
				   dir.c fat12.c fatreq.c open.c support.c \
				   names.c convers.c utf8.c utf16.c cp437.c \
				   case.c
	
	compile        -library=libextras.a fatinit.c
	
    cdl_option CYGPKG_FS_JFFS2_CFLAGS_ADD {
	display "Additional compiler flags"
	flavor  data
	no_define
	# We add -D__ECOS to trigger eCos-specific code in places.
	# We add -Werror because I find it useful.
	default_value { "-D__ECOS -nostdinc -iwithprefix include -Werror" }
	description   "
	    This option modifies the set of compiler flags for
            building the JFFS2 package.
            These flags are used in addition
            to the set of global flags."
        }

    cdl_option CYGPKG_FS_JFFS2_CFLAGS_REMOVE {
	display "Suppressed compiler flags"
	flavor  data
	no_define
	# We remove -Wpointer-arith so that some of the hacky Linux-compat code 
	# (in file.c) compiled. We can probably remove it when that's replaced
	# properly.
	default_value { "-Wpointer-arith" }
	description   "
	    This option modifies the set of compiler flags for
            building the JFFS2 package. These flags are removed from
            the set of global flags if present."
        }

    # ----------------------------------------------------------------
    # Tests

    cdl_option CYGPKG_FS_FAT_TESTS {
	display "FAT FS tests"
	flavor  data
	no_define
	calculated { "tests/fileio1" }
            description   "
                This option specifies the set of tests for the FAT FS package."
        }
    
}

# End of fat.cdl





