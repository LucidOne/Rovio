# ====================================================================
#
#      setjmp.cdl
#
#      C library setjmp/longjmp related configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jlarmour
# Contributors:
# Date:           2000-04-14
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_LIBC_SETJMP {
    display       "ISO C library setjmp/longjmp functions"
    description   "
        This package provides non-local jumps based on setjmp() and
        longjmp() in <setjmp.h> as specified by the ISO C
        standard - ISO/IEC 9899:1990."
    doc           ref/libc.html
    include_dir   cyg/libc/setjmp
    parent        CYGPKG_LIBC
    requires      CYGPKG_ISOINFRA
    implements    CYGINT_ISO_SETJMP
    requires      { CYGBLD_ISO_SETJMP_HEADER == "<cyg/libc/setjmp/setjmp.h>" }

    compile       longjmp.cxx

# ====================================================================


# ====================================================================

    cdl_component CYGPKG_LIBC_SETJMP_OPTIONS {
        display       "C library setjmp build options"
        flavor        none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_LIBC_SETJMP_CFLAGS_ADD {
            display       "Additional compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_LIBC_SETJMP_CFLAGS_REMOVE {
            display       "Suppressed compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_LIBC_SETJMP_TESTS {
            display       "C library setjmp tests"
            flavor        data
            no_define
            calculated    { "tests/setjmp" }
            description   "
                This option specifies the set of tests for this package."
        }
    }
}

# ====================================================================
# EOF setjmp.cdl
