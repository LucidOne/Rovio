# ====================================================================
#
#      termios.cdl
#
#      eCos POSIX termios compatible terminal configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jlarmour, gthomas
# Contributors:   
# Date:           2000-07-22
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_interface CYGINT_IO_SERIAL_TERMIOS_TERMIOS_TTY {
    display    "Interface for termios tty driver file enabling"
}

cdl_option CYGBLD_IO_SERIAL_TERMIOS_TERMIOS_TTY {
    display    "Build termios tty driver file"
    calculated 1
    active_if  { CYGINT_IO_SERIAL_TERMIOS_TERMIOS_TTY > 0 }
    compile    -library=libextras.a common/termiostty.c
}


cdl_component CYGPKG_IO_SERIAL_TERMIOS_TERMIOS0 {
    display       "Termios TTY channel #0"
    flavor        bool
    default_value 0
    implements    CYGINT_IO_SERIAL_TERMIOS_TERMIOS_TTY
    description   "
        This option causes '/dev/termios0' to be included in the standard 
        drivers."

    cdl_option CYGDAT_IO_SERIAL_TERMIOS_TERMIOS0_DEV {
        display       "Termios TTY channel #0 device"
        flavor        data
        default_value { "\"/dev/ser0\"" }
        description   "
            This option selects the physical device to use for 
            '/dev/termios0'."
    }
}
cdl_component CYGPKG_IO_SERIAL_TERMIOS_TERMIOS1 {
    display       "Termios TTY channel #1"
    flavor        bool
    default_value 0
    implements    CYGINT_IO_SERIAL_TERMIOS_TERMIOS_TTY
    description   "
        This option causes '/dev/termios1' to be included in the standard 
        drivers."

    cdl_option CYGDAT_IO_SERIAL_TERMIOS_TERMIOS1_DEV {
        display       "Termios TTY channel #1 device"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option selects the physical device to use for 
            '/dev/termios1'."
    }
}

cdl_component CYGPKG_IO_SERIAL_TERMIOS_TERMIOS2 {
    display       "Termios TTY channel #2"
    flavor        bool
    default_value 0
    implements    CYGINT_IO_SERIAL_TERMIOS_TERMIOS_TTY
    description   "
        This option causes '/dev/termios2' to be included in the standard 
        drivers."

    cdl_option CYGDAT_IO_SERIAL_TERMIOS_TERMIOS2_DEV {
        display       "Termios TTY channel #2 device"
        flavor        data
        default_value {"\"/dev/ser2\""}
        description   "
            This option selects the physical device to use for 
            '/dev/termios2'."
    }
}

cdl_option CYGSEM_IO_SERIAL_TERMIOS_USE_SIGNALS {
    display         "Support signals"
    flavor          bool
    requires        CYGINT_ISO_SIGNAL_NUMBERS
    requires        CYGINT_ISO_SIGNAL_IMPL
    default_value   { CYGINT_ISO_SIGNAL_NUMBERS != 0 && \
                      CYGINT_ISO_SIGNAL_IMPL != 0 }
    description     "This option selects whether those parts of the termios
                     interface involving signals is supported. This includes
                     BRKINT mode, the INTR and QUIT characters, and whether
                     SIGHUP is sent on terminal close."
}

# EOF termios.cdl
