# ====================================================================
#
#      bluetoothhci.cdl
#
#      bluetooth hci IO configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2004 Winbond.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      clyu
# Original data:  clyu
# Contributors:
# Date:           2004-08-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_BLUETOOTH_HCI {
    display       "Bluetooth HCI IO drivers"
    include_dir   cyg/io
    description   "
        This option enables drivers for basic I/O services on
        W99685 devices."
  	
  	requires       CYGPKG_LINUX_COMPAT
  	
    compile       -library=libextras.a	init.cxx hci_ldisc.c hci_h4.c

	 cdl_option CONFIG_BLUEZ_HCIUART_H4 {
        display		"blutooth hci uart h4 support"
        flavor        	bool
        default_value 	1
        description	"blutooth hci uart h4 support"
    }
    cdl_component CYGPKG_IO_BLUETOOTH_HCI_OPTIONS {
        display "Common W99685 support build options"
        flavor  none
		no_define

        cdl_option CYGPKG_IO_BLUETOOTH_HCI_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the common ethernet support package. These flags are used in addition
                to the set of global flags."
        }
    }
}
